  module test1;
     initial begin $display("Hello World"); $finish; end
  endmodule


